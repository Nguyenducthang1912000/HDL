library verilog;
use verilog.vl_types.all;
entity DMEM_vlg_check_tst is
    port(
        DATA_OUT        : in     vl_logic_vector(15 downto 0);
        sampler_rx      : in     vl_logic
    );
end DMEM_vlg_check_tst;
