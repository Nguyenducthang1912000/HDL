library verilog;
use verilog.vl_types.all;
entity AddConst_vlg_vec_tst is
end AddConst_vlg_vec_tst;
