library verilog;
use verilog.vl_types.all;
entity TestRF is
end TestRF;
