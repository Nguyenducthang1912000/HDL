library verilog;
use verilog.vl_types.all;
entity Inc2_vlg_vec_tst is
end Inc2_vlg_vec_tst;
