library verilog;
use verilog.vl_types.all;
entity TestStack is
end TestStack;
