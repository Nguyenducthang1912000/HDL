module 16bit_Processer (CLK);
//wire connection 
wire	PCSrc;
endmodule