library verilog;
use verilog.vl_types.all;
entity Cong_vlg_vec_tst is
end Cong_vlg_vec_tst;
