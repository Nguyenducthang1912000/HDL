library verilog;
use verilog.vl_types.all;
entity Lab1_vlg_check_tst is
    port(
        count_o         : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end Lab1_vlg_check_tst;
