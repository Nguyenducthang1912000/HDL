library verilog;
use verilog.vl_types.all;
entity Test_stack is
end Test_stack;
