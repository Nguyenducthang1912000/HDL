library verilog;
use verilog.vl_types.all;
entity Processer_16bit_vlg_vec_tst is
end Processer_16bit_vlg_vec_tst;
