library verilog;
use verilog.vl_types.all;
entity MooreFSM_vlg_vec_tst is
end MooreFSM_vlg_vec_tst;
