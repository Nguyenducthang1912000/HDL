library verilog;
use verilog.vl_types.all;
entity ASIC_vlg_vec_tst is
end ASIC_vlg_vec_tst;
