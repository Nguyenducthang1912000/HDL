library verilog;
use verilog.vl_types.all;
entity DMEM_vlg_vec_tst is
end DMEM_vlg_vec_tst;
