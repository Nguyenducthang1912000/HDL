library verilog;
use verilog.vl_types.all;
entity Processer_16bit_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Processer_16bit_vlg_sample_tst;
