library verilog;
use verilog.vl_types.all;
entity ShiftLeft1_vlg_vec_tst is
end ShiftLeft1_vlg_vec_tst;
